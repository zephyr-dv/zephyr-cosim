/****************************************************************************
 * zephyr_cosim.sv
 * 
 * Package provides SystemVerilog interface to Zephyr-Cosim
 ****************************************************************************/
  
/**
 * Package: zephyr_cosim
 * 
 * TODO: Add package documentation
 */
package zephyr_cosim;
	import tblink_rpc::*;

	class ZephyrCosim;
		
		function new();
		endfunction
		
		
	endclass


endpackage


