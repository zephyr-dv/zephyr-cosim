/****************************************************************************
 * sv_smoke_tb.sv
 ****************************************************************************/

/**
 * Module: sv_smoke_tb
 * 
 * TODO: Add module documentation
 */
module sv_smoke_tb(input clock);


endmodule


